module DELAY (input clk, input rst, output reg sig ,output reg err, output reg flg);
  localparam N = 200000;
  localparam CBITS = 18;
  reg [CBITS-1 :0] cnt;
  assign sig = (cnt >= N);
  assign err = (cnt > N);
  assign flg = (cnt < N);
  always @(posedge clk) begin
    if (rst || cnt >= N) cnt <= 0;
    else cnt <= cnt + 1; 
  end
	p1: assert property  ((@(posedge clk) sig |=> !sig)) ;
endmodule